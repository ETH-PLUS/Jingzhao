`timescale 1ns / 100ps
module cell_buf (
    input   A,
    output  Y
);

assign Y = A;

endmodule
