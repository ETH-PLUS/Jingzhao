module cell_clk_buf (
    input   A,
    output  Y
);

assign Y = A;

endmodule
