`ifndef HW_FORMAT_SV
`define HW_FORMAT_SV

`include "msg_def_v2p_h.vh"
`include "msg_def_ctxmgt_h.vh"
`include "ib_constant_def_h.vh"
`include "nic_hw_params.vh"
`include "sw_hw_interface_const_def_h.vh"

`define UNCERTAIN 0

`endif 
