`define SIMULATION
`define XILINX_FPGA
`define PCIEI_SIM
`define FPGA_VERSION

`define TD
