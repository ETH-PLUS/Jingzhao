//`define TD  #0.1
`define SIMPLE_MEM
`define FPGA_VERSION

//`define FPGA_V7_VALIDATE

`define VENDER_ID 16'h10EE
`define CAP_DSN   64'hA35_00000001

`define TD

`define XILINX_FPGA

`define ILA_ON

//`define ILA_HEADER_PARSER_ON
//`define ILA_PACKET_ENCAP_ON
//`define ILA_EXECUTION_ENGINE_ON
//`define ILA_VTP_ON
//`define ILA_CEU_ON
